module conventionToRBR(din, doutp, doutn);
	parameter no_of_digits = 8;
	input[no_of_digits-1:0] din;
	output[no_of_digits-1:0] doutp,doutn;
	
	

endmodule